-- Copyright (C) 1991-2011 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

library ieee;
use ieee.std_logic_1164.all;
library altera;
use altera.altera_syn_attributes.all;

entity reg_des is
	port
	(
		ck : in std_logic;
		d1 : in std_logic_vector(3 downto 0);
		d2 : in std_logic_vector(3 downto 0);
		ld : in std_logic;
		q1 : out std_logic_vector(3 downto 0);
		q2 : out std_logic_vector(3 downto 0)
	);

end reg_des;

architecture ppl_type of reg_des is

begin

end;
